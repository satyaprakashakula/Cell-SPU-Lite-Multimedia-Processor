module SPU_Lite_tb();
	
	logic clk, reset;
	//logic [0:7] IMem [1023:0];
	//logic [0:7] IMem_temp [1023:0];

	SPU_Lite SPU_Lite_inst(clk, reset);

	initial clk = 1;
	always #5 clk = ~clk;


	initial begin

		@(posedge clk); 
		#1; reset = 1; 

		/*
		IMem_temp [39:0] = '{
		'{8'b00011000}, '{8'b00001010}, '{8'b00001111}, '{8'b00010100}, 		  '{8'b00110001}, '{8'b00000000}, '{8'b00000101}, '{8'b00110010},  
		'{8'b00011000}, '{8'b00000000}, '{8'b11000001}, '{8'b00000001},           '{8'b00111011}, '{8'b01101000}, '{8'b00001111}, '{8'b10011110}, 
		'{8'b00011000}, '{8'b00000001}, '{8'b10000000}, '{8'b10000100},           '{8'b00111011}, '{8'b01101000}, '{8'b11000010}, '{8'b00100001}, 
		'{8'b00011000}, '{8'b00000010}, '{8'b01000100}, '{8'b00000111},			  '{8'b00111011}, '{8'b01101001}, '{8'b10010010}, '{8'b10100100}, 
		'{8'b00011000}, '{8'b00000010}, '{8'b10000101}, '{8'b10001100},           '{8'b00000000}, '{8'b00000000}, '{8'b00000000}, '{8'b00000000}
		};
		
		for(int i=0; i<40;i++) begin
			IMem[i] = IMem_temp[39-i]; 
		end

		for (int i=40; i<1024; i++) begin
			IMem[i] = 7'b0;
		end
		
		*/

		@(posedge clk); 
		#1; reset = 0;
		


		for(int i=0; i<300; i++) begin
			@(posedge clk);
		end


		$stop;


	end


endmodule






